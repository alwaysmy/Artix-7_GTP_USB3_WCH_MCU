module xillyusb_core
  (
  input  bus_clk,
  input  frontend_rst,
  input [31:0] pipe_rx,
  input  pipe_rx_clk,
  input [3:0] pipe_rx_k,
  input  pipe_rx_valid,
  input  pipe_tx_ready,
  input  pll_locked,
  input  receiver_present,
  input  receiver_present_valid,
  input  refclk_locked,
  input  rx_detect_revpolarity_clear,
  input  rx_elecidle,
  input  rx_phy_ready,
  input [7:0] user_r_mem_8_data,
  input  user_r_mem_8_empty,
  input  user_r_mem_8_eof,
  input [31:0] user_r_read_32_data,
  input  user_r_read_32_empty,
  input  user_r_read_32_eof,
  input [7:0] user_r_read_8_data,
  input  user_r_read_8_empty,
  input  user_r_read_8_eof,
  input  user_w_mem_8_full,
  input  user_w_write_32_full,
  input  user_w_write_8_full,
  input  version_gtp_1_0,
  output [7:0] gpio_led,
  output  lfps_en,
  output  mgt_en,
  output  mgt_powerdown,
  output [31:0] pipe_tx,
  output [3:0] pipe_tx_k,
  output  quiesce,
  output  receiver_detect,
  output  rx_align_enable,
  output  rx_detect_revpolarity,
  output  rx_dontmess,
  output  rx_resync,
  output [4:0] user_mem_8_addr,
  output  user_mem_8_addr_update,
  output  user_r_mem_8_open,
  output  user_r_mem_8_rden,
  output  user_r_read_32_open,
  output  user_r_read_32_rden,
  output  user_r_read_8_open,
  output  user_r_read_8_rden,
  output [7:0] user_w_mem_8_data,
  output  user_w_mem_8_open,
  output  user_w_mem_8_wren,
  output [31:0] user_w_write_32_data,
  output  user_w_write_32_open,
  output  user_w_write_32_wren,
  output [7:0] user_w_write_8_data,
  output  user_w_write_8_open,
  output  user_w_write_8_wren
);
endmodule
